library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;


entity main_mem is
    port (-- data buses
          addr         : in std_logic_vector(31 downto 0); 
          write_data   : in std_logic_vector(31 downto 0);
          read_data    : out std_logic_vector(31 downto 0);
          -- control signals
          Pet          : in std_logic;
          ReadOrWrite  : in std_logic;
          Ready        : out std_logic);
end data;

architecture Structure of main_mem is
    type ARRAY_MEM is array (2**8-1 downto 0) of std_logic_vector(7 downto 0);
    signal main_mem : ARRAY_MEM;
begin
    
    read_main_memory : process(Pet)
    begin
        if (Pet == '1' and ReadOrWrite == '0') then
            read_data(7 downto 0)    <= main_mem(to_integer(unsigned(addr      )));
            read_data(15 downto 8)   <= main_mem(to_integer(unsigned(addr+x"01")));
            read_data(23 downto 16)  <= main_mem(to_integer(unsigned(addr+x"02")));
            read_data(31 downto 24)  <= main_mem(to_integer(unsigned(addr+x"03")));
        end if;
        Ready <= '1';
    end process read_main_memory;

    write_main_memory : process(Pet)
    begin
        if (Pet == '1' and ReadOrWrite == '1') then
            main_mem(to_integer(unsigned(addr      ))) <= write_data(7 downto 0);
            main_mem(to_integer(unsigned(addr+x"01"))) <= write_data(15 downto 8);
            main_mem(to_integer(unsigned(addr+x"02"))) <= write_data(23 downto 16);
            main_mem(to_integer(unsigned(addr+x"03"))) <= write_data(31 downto 24); 
        end if;
        Ready <= '1';
    end process read_write_tags;

end Structure;
